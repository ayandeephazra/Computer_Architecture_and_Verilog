module seqdec_52(Inp, Clk, Reset, Out);
input Inp, Clk, Reset;
output Out;
wire reg1, reg2, reg3, reg4, reg5, reg6, reg7, reg8;
wire and1, and2, and3, and4, and5, and6, and7, and8;
dff iDFF1 (.q(reg1), .d(Inp), .clk(Clk), .rst(Reset));
dff iDFF2 (.q(reg2), .d(reg1), .clk(Clk), .rst(Reset));
dff iDFF3 (.q(reg3), .d(reg2), .clk(Clk), .rst(Reset));
dff iDFF4 (.q(reg4), .d(reg3), .clk(Clk), .rst(Reset));
dff iDFF5 (.q(reg5), .d(reg4), .clk(Clk), .rst(Reset));
dff iDFF6 (.q(reg6), .d(reg5), .clk(Clk), .rst(Reset));
dff iDFF7 (.q(reg7), .d(reg6), .clk(Clk), .rst(Reset));
dff iDFF8 (.q(reg8), .d(reg7), .clk(Clk), .rst(Reset));
not1 iNOT1(.in1(reg1), .out(and1));
assign and2 = reg2;
not1 iNOT2(.in1(reg3), .out(and3));
not1 iNOT3(.in1(reg4), .out(and4));
assign and5 = reg5;
not1 iNOT4(.in1(reg6), .out(and6));
assign and7 = reg7;
not1 iNOT5(.in1(reg8), .out(and8));

wire temp1, temp2, temp3, temp4, temp5, temp6, temp7, temp8, temp9, temp10, temp11, temp12, temp13, temp14;
nand2 iNAND2(.in1(and1),.in2(and2),.out(temp1));
not1 iNOT6(.in1(temp1), .out(temp2));
nand2 iNAND3(.in1(and3),.in2(temp2),.out(temp3));
not1 iNOT7(.in1(temp3), .out(temp4));
nand2 iNAND4(.in1(and4),.in2(temp4),.out(temp5));
not1 iNOT8(.in1(temp5), .out(temp6));
nand2 iNAND5(.in1(and5),.in2(temp6),.out(temp7));
not1 iNOT9(.in1(temp7), .out(temp8));
nand2 iNAND6(.in1(and6),.in2(temp8),.out(temp9));
not1 iNOT10(.in1(temp9), .out(temp10));
nand2 iNAND7(.in1(and7),.in2(temp10),.out(temp11));
not1 iNOT11(.in1(temp11), .out(temp12));
nand2 iNAND8(.in1(and8),.in2(temp12),.out(temp13));
not1 iNOT12(.in1(temp13), .out(temp14));
assign Out = temp14;
endmodule
