module proc_beqz_added (clk, rst, err);
    input clk;
    input rst;
    output err;

    // Your code

endmodule
