module branch_sel (op, zero, pos, neg, en);

  input [4:0] op;
  input zero, pos, neg;
  output reg en;

  always @(*) begin
    case (op)
///////////////////////////////////////////////////////////
// 		  	BEQZ		      		 // 
/////////////////////////////////////////////////////////// 
      5'b01100: en = (zero) ? 1'b1 : 1'b0;


///////////////////////////////////////////////////////////
// 		  	BNEZ		      		 // 
/////////////////////////////////////////////////////////// 
      5'b01101: en = (pos | neg) ? 1'b1 : 1'b0;


///////////////////////////////////////////////////////////
// 		  	BLTZ		      		 // 
/////////////////////////////////////////////////////////// 
      5'b01110: en = (neg) ? 1'b1 : 1'b0;


///////////////////////////////////////////////////////////
// 		  	BGEZ		      		 // 
/////////////////////////////////////////////////////////// 
      5'b01111: en = (pos | zero) ? 1'b1 : 1'b0;
      
      default: en = 1'b0;
    endcase

  end

endmodule