module fetch (clk, rst, beq_imm, err, instr);

	input clk;
	input rst;
	input [15:0] beq_imm;
	output err;
	output [15:0] instr;

	// Your Code goes here
	//reg [15:0] pc, pcPrev;
	wire [15:0] pcPrev_w;
	reg [15:0] A,B;
	
	wire[15:0] S, pc;
	wire Cout1, Cout2;
        wire [15:0] pc_fetch;
	wire [15:0] pc_u;
	wire [15:0] pc_beqmod;
////////////////////////////////
	memory2c iMEM(.data_out(instr), .data_in(16'h0000), .addr(pc_fetch), .enable(1'b1), .wr(1'b0), .createdump(1'b0), .clk(clk), .rst(rst));
	fulladder16 iFULLADDER1(.A(pc_fetch),.B(16'h0002),.S(pc_u),.Cout(Cout1));	
	fulladder16 iFULLADDER2(.A(pc_u),.B(beq_imm),.S(pc_beqmod),.Cout());	
        assign pc = (rst)? 16'h0000: pc_beqmod;
	dff IDFF [15:0] (.q(pc_fetch), .d(pc), .clk(clk), .rst(rst));


endmodule
