module fetch (clk, rst, err, instr);

	input clk;
	input rst;
	output err;
	output [15:0] instr;

	// Your Code goes here

endmodule
