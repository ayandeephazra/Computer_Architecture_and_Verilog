module control(instr, srcALU, regDestination, memWrite, regWrite, memtoreg, inv_A, inv_B, cin, AB, se, halt, siic, rti);

  input [15:0] instr;
  output reg [1:0] srcALU;
  output reg [1:0] regDestination;
  output reg memWrite, regWrite, memtoreg;
  output reg inv_A, inv_B, cin;
  output reg [4:0] AB;
  output reg se;
  output reg halt;
  output siic;
  output rti;

  assign siic = (instr[15:11]===5'b00010)? 1'b1: 1'b0;
  assign rti = (instr[15:11]===5'b00011)? 1'b1: 1'b0;  

  always @(*) begin
///////////////////////////////////////////////////////////////
// 	 	 DEFAULTING THE CONTROL SIGNALS  	     //
//	- - - - - - - - - - - - - - - - - - - - - - - -      //
//		memWrite, RegWrite, memtoreg -> 0	     //
//		       srcALU -> 0  			     //
//	   	       RegDst -> R7			     //
//			AB -> 0  			     //
//		inv_A, inv_B, Cin, se, halt -> 0	     //
///////////////////////////////////////////////////////////////
    srcALU = 2'b11; 
    regDestination = 2'b11; 
    memWrite = 1'b0;
    regWrite = 1'b0;
    memtoreg = 1'b0;
    inv_A = 1'b0;
    inv_B = 1'b0;
    cin = 1'b0;
    AB = 5'b00000;
    se = 1'b0;
    halt = 1'b0;
    //siic = 1'b0;
    //rti = 1'b0;

    case ({instr[15:11]})
///////////////////////////////////////////////////////////
// 		        HALT 		      		 //
//   Cease instruction issue, dump memory state to file	 //
/////////////////////////////////////////  //////////////// 
      5'b00000: begin 
        regDestination = 2'b00; 
        halt = 1'b1;
      end

///////////////////////////////////////////////////////////
// 		        NOP 		      		 //
//   			None				 //
/////////////////////////////////////////////////////////// 
      5'b00001: begin 
        regDestination = 2'b00; 
      end

///////////////////////////////////////////////////////////
// 		        ADDI 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b01000: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        AB = 5'b00010;
        se = 1'b1;
      end

///////////////////////////////////////////////////////////
// 		        SUBI 		      		 //
//   		    Rd, Rs, immediate			 //
///////////////////////////////////////////////////////////
      5'b01001: begin
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        inv_A = 1'b1;
        cin = 1'b1;
        AB = 5'b00010;
        se = 1'b1;
      end

///////////////////////////////////////////////////////////
// 		        XORI 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b01010: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        AB = 5'b00010;
      end

///////////////////////////////////////////////////////////
// 		        ANDI 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b01011: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        inv_B = 1'b1;
        AB = 5'b00010;
      end

///////////////////////////////////////////////////////////
// 		        ROLI 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10100: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        AB = 5'b00010;
      end

///////////////////////////////////////////////////////////
// 		        SLLI 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10101: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        AB = 5'b00010;
      end

///////////////////////////////////////////////////////////
// 		        RORI 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10110: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        AB = 5'b00010;
      end


///////////////////////////////////////////////////////////
// 		        SRLI 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10111: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        AB = 5'b00010;
      end

///////////////////////////////////////////////////////////
// 		        ST 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10000: begin 
        srcALU = 2'b01; 
        regDestination = 2'b10; 
        memWrite = 1'b1;
        AB = 5'b00011;
        se = 1'b1;
      end


///////////////////////////////////////////////////////////
// 		        LD 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10001: begin 
        srcALU = 2'b01; 
        regDestination = 2'b01; 
        regWrite = 1'b1;
        memtoreg = 1'b1;
        AB = 5'b00010;
        se = 1'b1;
      end


///////////////////////////////////////////////////////////
// 		        STU 		      		 //
//   		    Rd, Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10011: begin 
        srcALU = 2'b01; 
        regDestination = 2'b10; 
        memWrite = 1'b1;
        regWrite = 1'b1;
        AB = 5'b00011;
        se = 1'b1;
      end


///////////////////////////////////////////////////////////
// 		        BTR 		      		 //
//   		      Rd, Rs				 //
///////////////////////////////////////////////////////////
      5'b11001: begin 
        srcALU = 2'b11; 
        regDestination = 2'b00;
        regWrite = 1'b1;
        AB = 5'b00010;
      end


///////////////////////////////////////////////////////////
// 		  ADD/SUB/XOR/ANDN 	      		 //
//   		      Rd, Rs, Rt			 //
///////////////////////////////////////////////////////////
      5'b11011: begin 
        srcALU = 2'b00; 
        regDestination = 2'b00; 
        regWrite = 1'b1;
        inv_A = (instr[1:0] == 2'b01) ? 1'b1 : 1'b0;
        inv_B = (instr[1:0] == 2'b11) ? 1'b1 : 1'b0;
        cin = (instr[1:0] == 2'b01) ? 1'b1 : 1'b0;
        AB = 5'b00011;
      end

///////////////////////////////////////////////////////////
// 		  ROL/SLL/ROR/SRL	      		 //
//   		      Rd, Rs, Rt			 //
/////////////////////////////////////////////////////////// 
      5'b11010: begin 
        srcALU = 2'b00; 
        regDestination = 2'b00; 
        regWrite = 1'b1;
        AB = 5'b00011;
      end

///////////////////////////////////////////////////////////
// 		 	  SEQ      			 //
//   		      Rd, Rs, Rt			 //
///////////////////////////////////////////////////////////
      5'b11100: begin 
        srcALU = 2'b00; 
        regDestination = 2'b00; 
        regWrite = 1'b1;
        inv_B = 1'b1;
        cin = 1'b1;
        AB = 5'b00011;
      end

///////////////////////////////////////////////////////////
// 		  	SLT      	 		 //
//   		      Rd, Rs, Rt			 //
///////////////////////////////////////////////////////////
      5'b11101: begin 
        srcALU = 2'b00; 
        regDestination = 2'b00; 
        regWrite = 1'b1;
        inv_B = 1'b1;
        cin = 1'b1;
        AB = 5'b00011;
      end

///////////////////////////////////////////////////////////
// 		  	SLE      			 //
//   		      Rd, Rs, Rt			 //
/////////////////////////////////////////////////////////// 
      5'b11110: begin 
        srcALU = 2'b00; 
        regDestination = 2'b00; 
        regWrite = 1'b1;
        inv_B = 1'b1;
        cin = 1'b1;
        AB = 5'b00011;
      end

///////////////////////////////////////////////////////////
// 		  	SCO		      		 //
//   		      Rd, Rs, Rt			 //
/////////////////////////////////////////////////////////// 
      5'b11111: begin 
        srcALU = 2'b00; 
        regDestination = 2'b00; 
        regWrite = 1'b1;
        AB = 5'b00011;
      end

///////////////////////////////////////////////////////////
// 		  	BEQZ		      		 //
//   		     Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b01100: begin 
        regDestination = 2'b10; 
        inv_B = 1'b1;
        cin = 1'b1;
        AB = 5'b10010;
      end

///////////////////////////////////////////////////////////
// 		  	BNEZ		      		 //
//   		     Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b01101: begin 
        regDestination = 2'b10; 
        inv_B = 1'b1;
        cin = 1'b1;
        AB = 5'b10010;
      end

///////////////////////////////////////////////////////////
// 		  	BLTZ		      		 //
//   		     Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b01110: begin
        regDestination = 2'b10; 
        inv_B = 1'b1;
        cin = 1'b1;
        AB = 5'b10010;
      end


///////////////////////////////////////////////////////////
// 		  	BGEZ		      		 //
//   		     Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b01111: begin 
        regDestination = 2'b10; 
        inv_B = 1'b1;
        cin = 1'b1;
        AB = 5'b10010;
      end

///////////////////////////////////////////////////////////
// 		  	LBI		      		 //
//   		     Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b11000: begin 
        srcALU = 2'b10;
        regDestination = 2'b10; 
        regWrite = 1'b1;
        AB = 5'b00010;
        se = 1'b1;
      end

///////////////////////////////////////////////////////////
// 		  	SLBI		      		 //
//   		     Rs, immediate			 //
/////////////////////////////////////////////////////////// 
      5'b10010: begin 
        srcALU = 2'b10; 
        regDestination = 2'b10;
        regWrite = 1'b1;
        AB = 5'b00010;
      end

///////////////////////////////////////////////////////////
// 		  	J		      		 // 
///////////////////////////////////////////////////////////
      5'b00100: begin 
        AB = 5'b01000;
      end

///////////////////////////////////////////////////////////
// 		  	JR		      		 // 
/////////////////////////////////////////////////////////// 
      5'b00101: begin 
        AB = 5'b01010;
      end

///////////////////////////////////////////////////////////
// 		  	JAL		      		 // 
/////////////////////////////////////////////////////////// 
      5'b00110: begin 
        regWrite = 1'b1;
        AB = 5'b00100;
      end

///////////////////////////////////////////////////////////
// 		  	JALR		      		 // 
/////////////////////////////////////////////////////////// 
      5'b00111: begin 
        regWrite = 1'b1;
        AB = 5'b00110;
      end

///////////////////////////////////////////////////////////
// 		  	siic		      		 // 
/////////////////////////////////////////////////////////// 
      5'b00010: begin 
        regWrite = 1'b0;
        //siic = 1'b1;
      end

///////////////////////////////////////////////////////////
// 		  	NOP/RTI		      		 // 
/////////////////////////////////////////////////////////// 
      5'b00011: begin
        regWrite = 1'b0;
        //rti = 1'b1;
      end
      default: begin
      end
    endcase
  end
endmodule