 module proc(clk, rst, err);
    input clk;
    input rst;
    output err;

    // Your Code Here
endmodule
